`ifndef CONSTANTS_VH
`define CONSTANTS_VH

/* Incstucts Template
 * |15-13|12-10|9-7|6-4|3-0|
 */

`define INSTRUCT_ADD

`endif